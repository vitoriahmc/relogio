-- Copyright (C) 2016  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition
-- Created on Thu Sep 27 19:18:26 2018

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Z : IN STD_LOGIC := '0';
        palavra : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (IncrementaUS,ComparaUSCom9,ZeraUS,IncrementaDS,ComparaDSCom6,IncrementaUM,ZeraDS,ZeraUM,ComparaUMCom10,IncrementaDM,ComparaDMCom6,ZeraDM,IncrementaUH,ComparaUHCom4,ComparaDHCom2,ZeraUH,ZeraDH,ComparaUHCom10,ZeraUH_2,IncrementaDH);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_palavra : STD_LOGIC_VECTOR(14 DOWNTO 0) := "000000000000000";
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Z,reg_palavra)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= IncrementaUS;
            reg_palavra <= "000000000000000";
            palavra <= "000000000000000";
        ELSE
            reg_palavra <= "000000000000000";
            palavra <= "000000000000000";
            CASE fstate IS
                WHEN IncrementaUS =>
                    reg_fstate <= ComparaUSCom9;

                    reg_palavra <= "000000001001000";
                WHEN ComparaUSCom9 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= IncrementaUS;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= ZeraUS;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaUSCom9;
                    END IF;

                    reg_palavra <= "100000000101000";
                WHEN ZeraUS =>
                    reg_fstate <= IncrementaDS;

                    reg_palavra <= "010000001101000";
                WHEN IncrementaDS =>
                    reg_fstate <= ComparaDSCom6;

                    reg_palavra <= "000000010001001";
                WHEN ComparaDSCom6 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= IncrementaUS;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= ZeraDS;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaDSCom6;
                    END IF;

                    reg_palavra <= "100000000011001";
                WHEN IncrementaUM =>
                    reg_fstate <= ComparaUMCom10;

                    reg_palavra <= "000000100001010";
                WHEN ZeraDS =>
                    reg_fstate <= IncrementaUM;

                    reg_palavra <= "010000010011001";
                WHEN ZeraUM =>
                    reg_fstate <= IncrementaDM;

                    reg_palavra <= "010000100000010";
                WHEN ComparaUMCom10 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= IncrementaUS;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= ZeraUM;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaUMCom10;
                    END IF;

                    reg_palavra <= "100000000000010";
                WHEN IncrementaDM =>
                    reg_fstate <= ComparaDMCom6;

                    reg_palavra <= "000001000001011";
                WHEN ComparaDMCom6 =>
                    IF ((Z = '1')) THEN
                        reg_fstate <= ZeraDM;
                    ELSIF (NOT((Z = '1'))) THEN
                        reg_fstate <= IncrementaUS;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaDMCom6;
                    END IF;

                    reg_palavra <= "100000000011011";
                WHEN ZeraDM =>
                    reg_fstate <= IncrementaUH;

                    reg_palavra <= "010001000011011";
                WHEN IncrementaUH =>
                    reg_fstate <= ComparaUHCom4;

                    reg_palavra <= "000010000001100";
                WHEN ComparaUHCom4 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= ComparaUHCom10;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= ComparaDHCom2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaUHCom4;
                    END IF;

                    reg_palavra <= "100000000100100";
                WHEN ComparaDHCom2 =>
                    IF ((Z = '1')) THEN
                        reg_fstate <= ZeraUH;
                    ELSIF (NOT((Z = '1'))) THEN
                        reg_fstate <= IncrementaUS;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaDHCom2;
                    END IF;

                    reg_palavra <= "100000000010101";
                WHEN ZeraUH =>
                    reg_fstate <= ZeraDH;

                    reg_palavra <= "010010000100100";
                WHEN ZeraDH =>
                    reg_fstate <= IncrementaUS;

                    reg_palavra <= "010100000010101";
                WHEN ComparaUHCom10 =>
                    IF ((Z = '1')) THEN
                        reg_fstate <= ZeraUH_2;
                    ELSIF (NOT((Z = '1'))) THEN
                        reg_fstate <= IncrementaUS;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ComparaUHCom10;
                    END IF;

                    reg_palavra <= "100000000000100";
                WHEN ZeraUH_2 =>
                    reg_fstate <= IncrementaDH;

                    reg_palavra <= "010010000100100";
                WHEN IncrementaDH =>
                    reg_fstate <= IncrementaUS;

                    reg_palavra <= "000100000001101";
                WHEN OTHERS => 
                    reg_palavra <= "XXXXXXXXXXXXXXX";
                    report "Reach undefined state";
            END CASE;
            palavra <= reg_palavra;
        END IF;
    END PROCESS;
END BEHAVIOR;
